-------------------------------------------------------------------------------
-- Synthesizable syncronous 8-bit in 9-bit out ROM.
-- Outputs the input multiplied by c7 (as a signed integer).
-- 
-- Based on code by M. Treseler available at:
-- http://mysite.ncnetwork.net/reszotzl/sync_rom.vhd
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_rom_c7 is
    generic (data_length : natural := 8;
             add_length  : natural := 8);

    port ( clk          : in  std_logic;
           address      : in  std_logic_vector(add_length-1 downto 0);
           data_out     : out std_logic_vector(data_length-1 downto 0)
       );
end sync_rom_c7;

architecture synth_c7 of sync_rom_c7 is ---------------------------------------------
    constant mem_size : natural := 2**add_length;
    type     mem_type is array (mem_size-1 downto 0) of
    std_logic_vector (data_length-1 downto 0);
    constant mem : mem_type := (
       0 => "000000000" ,
       1 => "000000001" ,
       2 => "000000010" ,
       3 => "000000011" ,
       4 => "000000100" ,
       5 => "000000100" ,
       6 => "000000101" ,
       7 => "000000110" ,
       8 => "000000111" ,
       9 => "000001000" ,
       10 => "000001001" ,
       11 => "000001010" ,
       12 => "000001011" ,
       13 => "000001011" ,
       14 => "000001100" ,
       15 => "000001101" ,
       16 => "000001110" ,
       17 => "000001111" ,
       18 => "000010000" ,
       19 => "000010001" ,
       20 => "000010010" ,
       21 => "000010010" ,
       22 => "000010011" ,
       23 => "000010100" ,
       24 => "000010101" ,
       25 => "000010110" ,
       26 => "000010111" ,
       27 => "000011000" ,
       28 => "000011001" ,
       29 => "000011001" ,
       30 => "000011010" ,
       31 => "000011011" ,
       32 => "000011100" ,
       33 => "000011101" ,
       34 => "000011110" ,
       35 => "000011111" ,
       36 => "000100000" ,
       37 => "000100001" ,
       38 => "000100001" ,
       39 => "000100010" ,
       40 => "000100011" ,
       41 => "000100100" ,
       42 => "000100101" ,
       43 => "000100110" ,
       44 => "000100111" ,
       45 => "000101000" ,
       46 => "000101000" ,
       47 => "000101001" ,
       48 => "000101010" ,
       49 => "000101011" ,
       50 => "000101100" ,
       51 => "000101101" ,
       52 => "000101110" ,
       53 => "000101111" ,
       54 => "000101111" ,
       55 => "000110000" ,
       56 => "000110001" ,
       57 => "000110010" ,
       58 => "000110011" ,
       59 => "000110100" ,
       60 => "000110101" ,
       61 => "000110110" ,
       62 => "000110110" ,
       63 => "000110111" ,
       64 => "000111000" ,
       65 => "000111001" ,
       66 => "000111010" ,
       67 => "000111011" ,
       68 => "000111100" ,
       69 => "000111101" ,
       70 => "000111101" ,
       71 => "000111110" ,
       72 => "000111111" ,
       73 => "001000000" ,
       74 => "001000001" ,
       75 => "001000010" ,
       76 => "001000011" ,
       77 => "001000100" ,
       78 => "001000101" ,
       79 => "001000101" ,
       80 => "001000110" ,
       81 => "001000111" ,
       82 => "001001000" ,
       83 => "001001001" ,
       84 => "001001010" ,
       85 => "001001011" ,
       86 => "001001100" ,
       87 => "001001100" ,
       88 => "001001101" ,
       89 => "001001110" ,
       90 => "001001111" ,
       91 => "001010000" ,
       92 => "001010001" ,
       93 => "001010010" ,
       94 => "001010011" ,
       95 => "001010011" ,
       96 => "001010100" ,
       97 => "001010101" ,
       98 => "001010110" ,
       99 => "001010111" ,
       100 => "001011000" ,
       101 => "001011001" ,
       102 => "001011010" ,
       103 => "001011010" ,
       104 => "001011011" ,
       105 => "001011100" ,
       106 => "001011101" ,
       107 => "001011110" ,
       108 => "001011111" ,
       109 => "001100000" ,
       110 => "001100001" ,
       111 => "001100010" ,
       112 => "001100010" ,
       113 => "001100011" ,
       114 => "001100100" ,
       115 => "001100101" ,
       116 => "001100110" ,
       117 => "001100111" ,
       118 => "001101000" ,
       119 => "001101001" ,
       120 => "001101001" ,
       121 => "001101010" ,
       122 => "001101011" ,
       123 => "001101100" ,
       124 => "001101101" ,
       125 => "001101110" ,
       126 => "001101111" ,
       127 => "001110000" ,
       128 => "001110000" ,
       129 => "001110001" ,
       130 => "001110010" ,
       131 => "001110011" ,
       132 => "001110100" ,
       133 => "001110101" ,
       134 => "001110110" ,
       135 => "001110111" ,
       136 => "001110111" ,
       137 => "001111000" ,
       138 => "001111001" ,
       139 => "001111010" ,
       140 => "001111011" ,
       141 => "001111100" ,
       142 => "001111101" ,
       143 => "001111110" ,
       144 => "001111110" ,
       145 => "001111111" ,
       146 => "010000000" ,
       147 => "010000001" ,
       148 => "010000010" ,
       149 => "010000011" ,
       150 => "010000100" ,
       151 => "010000101" ,
       152 => "010000110" ,
       153 => "010000110" ,
       154 => "010000111" ,
       155 => "010001000" ,
       156 => "010001001" ,
       157 => "010001010" ,
       158 => "010001011" ,
       159 => "010001100" ,
       160 => "010001101" ,
       161 => "010001101" ,
       162 => "010001110" ,
       163 => "010001111" ,
       164 => "010010000" ,
       165 => "010010001" ,
       166 => "010010010" ,
       167 => "010010011" ,
       168 => "010010100" ,
       169 => "010010100" ,
       170 => "010010101" ,
       171 => "010010110" ,
       172 => "010010111" ,
       173 => "010011000" ,
       174 => "010011001" ,
       175 => "010011010" ,
       176 => "010011011" ,
       177 => "010011011" ,
       178 => "010011100" ,
       179 => "010011101" ,
       180 => "010011110" ,
       181 => "010011111" ,
       182 => "010100000" ,
       183 => "010100001" ,
       184 => "010100010" ,
       185 => "010100011" ,
       186 => "010100011" ,
       187 => "010100100" ,
       188 => "010100101" ,
       189 => "010100110" ,
       190 => "010100111" ,
       191 => "010101000" ,
       192 => "010101001" ,
       193 => "010101010" ,
       194 => "010101010" ,
       195 => "010101011" ,
       196 => "010101100" ,
       197 => "010101101" ,
       198 => "010101110" ,
       199 => "010101111" ,
       200 => "010110000" ,
       201 => "010110001" ,
       202 => "010110001" ,
       203 => "010110010" ,
       204 => "010110011" ,
       205 => "010110100" ,
       206 => "010110101" ,
       207 => "010110110" ,
       208 => "010110111" ,
       209 => "010111000" ,
       210 => "010111000" ,
       211 => "010111001" ,
       212 => "010111010" ,
       213 => "010111011" ,
       214 => "010111100" ,
       215 => "010111101" ,
       216 => "010111110" ,
       217 => "010111111" ,
       218 => "010111111" ,
       219 => "011000000" ,
       220 => "011000001" ,
       221 => "011000010" ,
       222 => "011000011" ,
       223 => "011000100" ,
       224 => "011000101" ,
       225 => "011000110" ,
       226 => "011000111" ,
       227 => "011000111" ,
       228 => "011001000" ,
       229 => "011001001" ,
       230 => "011001010" ,
       231 => "011001011" ,
       232 => "011001100" ,
       233 => "011001101" ,
       234 => "011001110" ,
       235 => "011001110" ,
       236 => "011001111" ,
       237 => "011010000" ,
       238 => "011010001" ,
       239 => "011010010" ,
       240 => "011010011" ,
       241 => "011010100" ,
       242 => "011010101" ,
       243 => "011010101" ,
       244 => "011010110" ,
       245 => "011010111" ,
       246 => "011011000" ,
       247 => "011011001" ,
       248 => "011011010" ,
       249 => "011011011" ,
       250 => "011011100" ,
       251 => "011011100" ,
       252 => "011011101" ,
       253 => "011011110" ,
       254 => "011011111" ,
       255 => "011100000"
    );

begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <= mem(to_integer(unsigned(address))); 
        end if;
    end process rom;

end architecture synth_c7;

