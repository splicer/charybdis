-------------------------------------------------------------------------------
-- Synthesizable syncronous 8-bit in 9-bit out ROM.
-- Outputs the input multiplied by c8 (as a signed integer).
-- 
-- Based on code by M. Treseler available at:
-- http://mysite.ncnetwork.net/reszotzl/sync_rom.vhd
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_rom_c8 is
    generic (data_length : natural := 9;
             add_length  : natural := 8);

    port ( clk          : in  std_logic;
           address      : in  std_logic_vector(add_length-1 downto 0);
           data_out     : out std_logic_vector(data_length-1 downto 0)
       );
end sync_rom_c8;

architecture synth_c8 of sync_rom_c8 is ---------------------------------------------
    constant mem_size : natural := 2**add_length;
    type     mem_type is array (mem_size-1 downto 0) of
    std_logic_vector (data_length-1 downto 0);
    constant mem : mem_type := (
       0 => "000000000" ,
       1 => "111111111" ,
       2 => "111111111" ,
       3 => "111111110" ,
       4 => "111111101" ,
       5 => "111111100" ,
       6 => "111111100" ,
       7 => "111111011" ,
       8 => "111111010" ,
       9 => "111111001" ,
       10 => "111111001" ,
       11 => "111111000" ,
       12 => "111110111" ,
       13 => "111110110" ,
       14 => "111110110" ,
       15 => "111110101" ,
       16 => "111110100" ,
       17 => "111110011" ,
       18 => "111110011" ,
       19 => "111110010" ,
       20 => "111110001" ,
       21 => "111110001" ,
       22 => "111110000" ,
       23 => "111101111" ,
       24 => "111101110" ,
       25 => "111101110" ,
       26 => "111101101" ,
       27 => "111101100" ,
       28 => "111101011" ,
       29 => "111101011" ,
       30 => "111101010" ,
       31 => "111101001" ,
       32 => "111101000" ,
       33 => "111101000" ,
       34 => "111100111" ,
       35 => "111100110" ,
       36 => "111100110" ,
       37 => "111100101" ,
       38 => "111100100" ,
       39 => "111100011" ,
       40 => "111100011" ,
       41 => "111100010" ,
       42 => "111100001" ,
       43 => "111100000" ,
       44 => "111100000" ,
       45 => "111011111" ,
       46 => "111011110" ,
       47 => "111011101" ,
       48 => "111011101" ,
       49 => "111011100" ,
       50 => "111011011" ,
       51 => "111011010" ,
       52 => "111011010" ,
       53 => "111011001" ,
       54 => "111011000" ,
       55 => "111011000" ,
       56 => "111010111" ,
       57 => "111010110" ,
       58 => "111010101" ,
       59 => "111010101" ,
       60 => "111010100" ,
       61 => "111010011" ,
       62 => "111010010" ,
       63 => "111010010" ,
       64 => "111010001" ,
       65 => "111010000" ,
       66 => "111001111" ,
       67 => "111001111" ,
       68 => "111001110" ,
       69 => "111001101" ,
       70 => "111001101" ,
       71 => "111001100" ,
       72 => "111001011" ,
       73 => "111001010" ,
       74 => "111001010" ,
       75 => "111001001" ,
       76 => "111001000" ,
       77 => "111000111" ,
       78 => "111000111" ,
       79 => "111000110" ,
       80 => "111000101" ,
       81 => "111000100" ,
       82 => "111000100" ,
       83 => "111000011" ,
       84 => "111000010" ,
       85 => "111000001" ,
       86 => "111000001" ,
       87 => "111000000" ,
       88 => "110111111" ,
       89 => "110111111" ,
       90 => "110111110" ,
       91 => "110111101" ,
       92 => "110111100" ,
       93 => "110111100" ,
       94 => "110111011" ,
       95 => "110111010" ,
       96 => "110111001" ,
       97 => "110111001" ,
       98 => "110111000" ,
       99 => "110110111" ,
       100 => "110110110" ,
       101 => "110110110" ,
       102 => "110110101" ,
       103 => "110110100" ,
       104 => "110110011" ,
       105 => "110110011" ,
       106 => "110110010" ,
       107 => "110110001" ,
       108 => "110110001" ,
       109 => "110110000" ,
       110 => "110101111" ,
       111 => "110101110" ,
       112 => "110101110" ,
       113 => "110101101" ,
       114 => "110101100" ,
       115 => "110101011" ,
       116 => "110101011" ,
       117 => "110101010" ,
       118 => "110101001" ,
       119 => "110101000" ,
       120 => "110101000" ,
       121 => "110100111" ,
       122 => "110100110" ,
       123 => "110100110" ,
       124 => "110100101" ,
       125 => "110100100" ,
       126 => "110100011" ,
       127 => "110100011" ,
       128 => "110100010" ,
       129 => "110100001" ,
       130 => "110100000" ,
       131 => "110100000" ,
       132 => "110011111" ,
       133 => "110011110" ,
       134 => "110011101" ,
       135 => "110011101" ,
       136 => "110011100" ,
       137 => "110011011" ,
       138 => "110011010" ,
       139 => "110011010" ,
       140 => "110011001" ,
       141 => "110011000" ,
       142 => "110011000" ,
       143 => "110010111" ,
       144 => "110010110" ,
       145 => "110010101" ,
       146 => "110010101" ,
       147 => "110010100" ,
       148 => "110010011" ,
       149 => "110010010" ,
       150 => "110010010" ,
       151 => "110010001" ,
       152 => "110010000" ,
       153 => "110001111" ,
       154 => "110001111" ,
       155 => "110001110" ,
       156 => "110001101" ,
       157 => "110001101" ,
       158 => "110001100" ,
       159 => "110001011" ,
       160 => "110001010" ,
       161 => "110001010" ,
       162 => "110001001" ,
       163 => "110001000" ,
       164 => "110000111" ,
       165 => "110000111" ,
       166 => "110000110" ,
       167 => "110000101" ,
       168 => "110000100" ,
       169 => "110000100" ,
       170 => "110000011" ,
       171 => "110000010" ,
       172 => "110000001" ,
       173 => "110000001" ,
       174 => "110000000" ,
       175 => "101111111" ,
       176 => "101111111" ,
       177 => "101111110" ,
       178 => "101111101" ,
       179 => "101111100" ,
       180 => "101111100" ,
       181 => "101111011" ,
       182 => "101111010" ,
       183 => "101111001" ,
       184 => "101111001" ,
       185 => "101111000" ,
       186 => "101110111" ,
       187 => "101110110" ,
       188 => "101110110" ,
       189 => "101110101" ,
       190 => "101110100" ,
       191 => "101110100" ,
       192 => "101110011" ,
       193 => "101110010" ,
       194 => "101110001" ,
       195 => "101110001" ,
       196 => "101110000" ,
       197 => "101101111" ,
       198 => "101101110" ,
       199 => "101101110" ,
       200 => "101101101" ,
       201 => "101101100" ,
       202 => "101101011" ,
       203 => "101101011" ,
       204 => "101101010" ,
       205 => "101101001" ,
       206 => "101101000" ,
       207 => "101101000" ,
       208 => "101100111" ,
       209 => "101100110" ,
       210 => "101100110" ,
       211 => "101100101" ,
       212 => "101100100" ,
       213 => "101100011" ,
       214 => "101100011" ,
       215 => "101100010" ,
       216 => "101100001" ,
       217 => "101100000" ,
       218 => "101100000" ,
       219 => "101011111" ,
       220 => "101011110" ,
       221 => "101011101" ,
       222 => "101011101" ,
       223 => "101011100" ,
       224 => "101011011" ,
       225 => "101011010" ,
       226 => "101011010" ,
       227 => "101011001" ,
       228 => "101011000" ,
       229 => "101011000" ,
       230 => "101010111" ,
       231 => "101010110" ,
       232 => "101010101" ,
       233 => "101010101" ,
       234 => "101010100" ,
       235 => "101010011" ,
       236 => "101010010" ,
       237 => "101010010" ,
       238 => "101010001" ,
       239 => "101010000" ,
       240 => "101001111" ,
       241 => "101001111" ,
       242 => "101001110" ,
       243 => "101001101" ,
       244 => "101001101" ,
       245 => "101001100" ,
       246 => "101001011" ,
       247 => "101001010" ,
       248 => "101001010" ,
       249 => "101001001" ,
       250 => "101001000" ,
       251 => "101000111" ,
       252 => "101000111" ,
       253 => "101000110" ,
       254 => "101000101" ,
       255 => "101000100"
    );

begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <= mem(to_integer(unsigned(address))); 
        end if;
    end process rom;

end architecture synth_c8;

