-------------------------------------------------------------------------------
-- Synthesizable syncronous 8-bit in 8-bit out ROM.
-- Outputs the input multiplied by c1 (as an unsigned integer).
-- 
-- Based on code by M. Treseler available at:
-- http://mysite.ncnetwork.net/reszotzl/sync_rom.vhd
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_rom_c1 is
    generic (data_length : natural := 8;
             add_length  : natural := 8);

    port ( clk          : in  std_logic;
           address      : in  std_logic_vector(add_length-1 downto 0);
           data_out     : out std_logic_vector(data_length-1 downto 0)
       );
end sync_rom_c1;

architecture synth_c1 of sync_rom_c1 is ---------------------------------------------
    constant mem_size : natural := 2**add_length;
    type     mem_type is array (mem_size-1 downto 0) of
    std_logic_vector (data_length-1 downto 0);
    constant mem : mem_type := (
        0 => "00000000" ,
        1 => "00000000" ,
        2 => "00000001" ,
        3 => "00000001" ,
        4 => "00000001" ,
        5 => "00000001" ,
        6 => "00000010" ,
        7 => "00000010" ,
        8 => "00000010" ,
        9 => "00000010" ,
        10 => "00000011" ,
        11 => "00000011" ,
        12 => "00000011" ,
        13 => "00000011" ,
        14 => "00000100" ,
        15 => "00000100" ,
        16 => "00000100" ,
        17 => "00000100" ,
        18 => "00000101" ,
        19 => "00000101" ,
        20 => "00000101" ,
        21 => "00000101" ,
        22 => "00000110" ,
        23 => "00000110" ,
        24 => "00000110" ,
        25 => "00000110" ,
        26 => "00000111" ,
        27 => "00000111" ,
        28 => "00000111" ,
        29 => "00000111" ,
        30 => "00001000" ,
        31 => "00001000" ,
        32 => "00001000" ,
        33 => "00001000" ,
        34 => "00001001" ,
        35 => "00001001" ,
        36 => "00001001" ,
        37 => "00001010" ,
        38 => "00001010" ,
        39 => "00001010" ,
        40 => "00001010" ,
        41 => "00001011" ,
        42 => "00001011" ,
        43 => "00001011" ,
        44 => "00001011" ,
        45 => "00001100" ,
        46 => "00001100" ,
        47 => "00001100" ,
        48 => "00001100" ,
        49 => "00001101" ,
        50 => "00001101" ,
        51 => "00001101" ,
        52 => "00001101" ,
        53 => "00001110" ,
        54 => "00001110" ,
        55 => "00001110" ,
        56 => "00001110" ,
        57 => "00001111" ,
        58 => "00001111" ,
        59 => "00001111" ,
        60 => "00001111" ,
        61 => "00010000" ,
        62 => "00010000" ,
        63 => "00010000" ,
        64 => "00010000" ,
        65 => "00010001" ,
        66 => "00010001" ,
        67 => "00010001" ,
        68 => "00010001" ,
        69 => "00010010" ,
        70 => "00010010" ,
        71 => "00010010" ,
        72 => "00010010" ,
        73 => "00010011" ,
        74 => "00010011" ,
        75 => "00010011" ,
        76 => "00010100" ,
        77 => "00010100" ,
        78 => "00010100" ,
        79 => "00010100" ,
        80 => "00010101" ,
        81 => "00010101" ,
        82 => "00010101" ,
        83 => "00010101" ,
        84 => "00010110" ,
        85 => "00010110" ,
        86 => "00010110" ,
        87 => "00010110" ,
        88 => "00010111" ,
        89 => "00010111" ,
        90 => "00010111" ,
        91 => "00010111" ,
        92 => "00011000" ,
        93 => "00011000" ,
        94 => "00011000" ,
        95 => "00011000" ,
        96 => "00011001" ,
        97 => "00011001" ,
        98 => "00011001" ,
        99 => "00011001" ,
        100 => "00011010" ,
        101 => "00011010" ,
        102 => "00011010" ,
        103 => "00011010" ,
        104 => "00011011" ,
        105 => "00011011" ,
        106 => "00011011" ,
        107 => "00011011" ,
        108 => "00011100" ,
        109 => "00011100" ,
        110 => "00011100" ,
        111 => "00011101" ,
        112 => "00011101" ,
        113 => "00011101" ,
        114 => "00011101" ,
        115 => "00011110" ,
        116 => "00011110" ,
        117 => "00011110" ,
        118 => "00011110" ,
        119 => "00011111" ,
        120 => "00011111" ,
        121 => "00011111" ,
        122 => "00011111" ,
        123 => "00100000" ,
        124 => "00100000" ,
        125 => "00100000" ,
        126 => "00100000" ,
        127 => "00100001" ,
        128 => "00100001" ,
        129 => "00100001" ,
        130 => "00100001" ,
        131 => "00100010" ,
        132 => "00100010" ,
        133 => "00100010" ,
        134 => "00100010" ,
        135 => "00100011" ,
        136 => "00100011" ,
        137 => "00100011" ,
        138 => "00100011" ,
        139 => "00100100" ,
        140 => "00100100" ,
        141 => "00100100" ,
        142 => "00100100" ,
        143 => "00100101" ,
        144 => "00100101" ,
        145 => "00100101" ,
        146 => "00100101" ,
        147 => "00100110" ,
        148 => "00100110" ,
        149 => "00100110" ,
        150 => "00100111" ,
        151 => "00100111" ,
        152 => "00100111" ,
        153 => "00100111" ,
        154 => "00101000" ,
        155 => "00101000" ,
        156 => "00101000" ,
        157 => "00101000" ,
        158 => "00101001" ,
        159 => "00101001" ,
        160 => "00101001" ,
        161 => "00101001" ,
        162 => "00101010" ,
        163 => "00101010" ,
        164 => "00101010" ,
        165 => "00101010" ,
        166 => "00101011" ,
        167 => "00101011" ,
        168 => "00101011" ,
        169 => "00101011" ,
        170 => "00101100" ,
        171 => "00101100" ,
        172 => "00101100" ,
        173 => "00101100" ,
        174 => "00101101" ,
        175 => "00101101" ,
        176 => "00101101" ,
        177 => "00101101" ,
        178 => "00101110" ,
        179 => "00101110" ,
        180 => "00101110" ,
        181 => "00101110" ,
        182 => "00101111" ,
        183 => "00101111" ,
        184 => "00101111" ,
        185 => "00110000" ,
        186 => "00110000" ,
        187 => "00110000" ,
        188 => "00110000" ,
        189 => "00110001" ,
        190 => "00110001" ,
        191 => "00110001" ,
        192 => "00110001" ,
        193 => "00110010" ,
        194 => "00110010" ,
        195 => "00110010" ,
        196 => "00110010" ,
        197 => "00110011" ,
        198 => "00110011" ,
        199 => "00110011" ,
        200 => "00110011" ,
        201 => "00110100" ,
        202 => "00110100" ,
        203 => "00110100" ,
        204 => "00110100" ,
        205 => "00110101" ,
        206 => "00110101" ,
        207 => "00110101" ,
        208 => "00110101" ,
        209 => "00110110" ,
        210 => "00110110" ,
        211 => "00110110" ,
        212 => "00110110" ,
        213 => "00110111" ,
        214 => "00110111" ,
        215 => "00110111" ,
        216 => "00110111" ,
        217 => "00111000" ,
        218 => "00111000" ,
        219 => "00111000" ,
        220 => "00111000" ,
        221 => "00111001" ,
        222 => "00111001" ,
        223 => "00111001" ,
        224 => "00111010" ,
        225 => "00111010" ,
        226 => "00111010" ,
        227 => "00111010" ,
        228 => "00111011" ,
        229 => "00111011" ,
        230 => "00111011" ,
        231 => "00111011" ,
        232 => "00111100" ,
        233 => "00111100" ,
        234 => "00111100" ,
        235 => "00111100" ,
        236 => "00111101" ,
        237 => "00111101" ,
        238 => "00111101" ,
        239 => "00111101" ,
        240 => "00111110" ,
        241 => "00111110" ,
        242 => "00111110" ,
        243 => "00111110" ,
        244 => "00111111" ,
        245 => "00111111" ,
        246 => "00111111" ,
        247 => "00111111" ,
        248 => "01000000" ,
        249 => "01000000" ,
        250 => "01000000" ,
        251 => "01000000" ,
        252 => "01000001" ,
        253 => "01000001" ,
        254 => "01000001" ,
        255 => "01000001"
    );

begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <= mem(to_integer(unsigned(address))); 
        end if;
    end process rom;

end architecture synth_c1;

