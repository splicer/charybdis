-------------------------------------------------------------------------------
-- Synthesizable syncronous 8-bit in 9-bit out ROM.
-- Outputs the input multiplied by c9 (as a signed integer).
-- 
-- Based on code by M. Treseler available at:
-- http://mysite.ncnetwork.net/reszotzl/sync_rom.vhd
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_rom_c9 is
    generic (data_length : natural := 9;
             add_length  : natural := 8);

    port ( clk          : in  std_logic;
           address      : in  std_logic_vector(add_length-1 downto 0);
           data_out     : out std_logic_vector(data_length-1 downto 0)
       );
end sync_rom_c9;

architecture synth_c9 of sync_rom_c9 is ---------------------------------------------
    constant mem_size : natural := 2**add_length;
    type     mem_type is array (mem_size-1 downto 0) of
    std_logic_vector (data_length-1 downto 0);
    constant mem : mem_type := (
        0 => "000000000" ,
        1 => "000000000" ,
        2 => "000000000" ,
        3 => "000000000" ,
        4 => "111111111" ,
        5 => "111111111" ,
        6 => "111111111" ,
        7 => "111111111" ,
        8 => "111111111" ,
        9 => "111111111" ,
        10 => "111111111" ,
        11 => "111111110" ,
        12 => "111111110" ,
        13 => "111111110" ,
        14 => "111111110" ,
        15 => "111111110" ,
        16 => "111111110" ,
        17 => "111111110" ,
        18 => "111111101" ,
        19 => "111111101" ,
        20 => "111111101" ,
        21 => "111111101" ,
        22 => "111111101" ,
        23 => "111111101" ,
        24 => "111111101" ,
        25 => "111111100" ,
        26 => "111111100" ,
        27 => "111111100" ,
        28 => "111111100" ,
        29 => "111111100" ,
        30 => "111111100" ,
        31 => "111111100" ,
        32 => "111111011" ,
        33 => "111111011" ,
        34 => "111111011" ,
        35 => "111111011" ,
        36 => "111111011" ,
        37 => "111111011" ,
        38 => "111111011" ,
        39 => "111111010" ,
        40 => "111111010" ,
        41 => "111111010" ,
        42 => "111111010" ,
        43 => "111111010" ,
        44 => "111111010" ,
        45 => "111111010" ,
        46 => "111111001" ,
        47 => "111111001" ,
        48 => "111111001" ,
        49 => "111111001" ,
        50 => "111111001" ,
        51 => "111111001" ,
        52 => "111111001" ,
        53 => "111111000" ,
        54 => "111111000" ,
        55 => "111111000" ,
        56 => "111111000" ,
        57 => "111111000" ,
        58 => "111111000" ,
        59 => "111111000" ,
        60 => "111110111" ,
        61 => "111110111" ,
        62 => "111110111" ,
        63 => "111110111" ,
        64 => "111110111" ,
        65 => "111110111" ,
        66 => "111110111" ,
        67 => "111110110" ,
        68 => "111110110" ,
        69 => "111110110" ,
        70 => "111110110" ,
        71 => "111110110" ,
        72 => "111110110" ,
        73 => "111110110" ,
        74 => "111110101" ,
        75 => "111110101" ,
        76 => "111110101" ,
        77 => "111110101" ,
        78 => "111110101" ,
        79 => "111110101" ,
        80 => "111110101" ,
        81 => "111110100" ,
        82 => "111110100" ,
        83 => "111110100" ,
        84 => "111110100" ,
        85 => "111110100" ,
        86 => "111110100" ,
        87 => "111110100" ,
        88 => "111110011" ,
        89 => "111110011" ,
        90 => "111110011" ,
        91 => "111110011" ,
        92 => "111110011" ,
        93 => "111110011" ,
        94 => "111110011" ,
        95 => "111110010" ,
        96 => "111110010" ,
        97 => "111110010" ,
        98 => "111110010" ,
        99 => "111110010" ,
        100 => "111110010" ,
        101 => "111110010" ,
        102 => "111110001" ,
        103 => "111110001" ,
        104 => "111110001" ,
        105 => "111110001" ,
        106 => "111110001" ,
        107 => "111110001" ,
        108 => "111110001" ,
        109 => "111110000" ,
        110 => "111110000" ,
        111 => "111110000" ,
        112 => "111110000" ,
        113 => "111110000" ,
        114 => "111110000" ,
        115 => "111110000" ,
        116 => "111101111" ,
        117 => "111101111" ,
        118 => "111101111" ,
        119 => "111101111" ,
        120 => "111101111" ,
        121 => "111101111" ,
        122 => "111101111" ,
        123 => "111101110" ,
        124 => "111101110" ,
        125 => "111101110" ,
        126 => "111101110" ,
        127 => "111101110" ,
        128 => "111101110" ,
        129 => "111101110" ,
        130 => "111101101" ,
        131 => "111101101" ,
        132 => "111101101" ,
        133 => "111101101" ,
        134 => "111101101" ,
        135 => "111101101" ,
        136 => "111101101" ,
        137 => "111101100" ,
        138 => "111101100" ,
        139 => "111101100" ,
        140 => "111101100" ,
        141 => "111101100" ,
        142 => "111101100" ,
        143 => "111101100" ,
        144 => "111101011" ,
        145 => "111101011" ,
        146 => "111101011" ,
        147 => "111101011" ,
        148 => "111101011" ,
        149 => "111101011" ,
        150 => "111101011" ,
        151 => "111101010" ,
        152 => "111101010" ,
        153 => "111101010" ,
        154 => "111101010" ,
        155 => "111101010" ,
        156 => "111101010" ,
        157 => "111101010" ,
        158 => "111101001" ,
        159 => "111101001" ,
        160 => "111101001" ,
        161 => "111101001" ,
        162 => "111101001" ,
        163 => "111101001" ,
        164 => "111101001" ,
        165 => "111101000" ,
        166 => "111101000" ,
        167 => "111101000" ,
        168 => "111101000" ,
        169 => "111101000" ,
        170 => "111101000" ,
        171 => "111101000" ,
        172 => "111100111" ,
        173 => "111100111" ,
        174 => "111100111" ,
        175 => "111100111" ,
        176 => "111100111" ,
        177 => "111100111" ,
        178 => "111100111" ,
        179 => "111100110" ,
        180 => "111100110" ,
        181 => "111100110" ,
        182 => "111100110" ,
        183 => "111100110" ,
        184 => "111100110" ,
        185 => "111100110" ,
        186 => "111100101" ,
        187 => "111100101" ,
        188 => "111100101" ,
        189 => "111100101" ,
        190 => "111100101" ,
        191 => "111100101" ,
        192 => "111100101" ,
        193 => "111100100" ,
        194 => "111100100" ,
        195 => "111100100" ,
        196 => "111100100" ,
        197 => "111100100" ,
        198 => "111100100" ,
        199 => "111100100" ,
        200 => "111100011" ,
        201 => "111100011" ,
        202 => "111100011" ,
        203 => "111100011" ,
        204 => "111100011" ,
        205 => "111100011" ,
        206 => "111100011" ,
        207 => "111100010" ,
        208 => "111100010" ,
        209 => "111100010" ,
        210 => "111100010" ,
        211 => "111100010" ,
        212 => "111100010" ,
        213 => "111100010" ,
        214 => "111100001" ,
        215 => "111100001" ,
        216 => "111100001" ,
        217 => "111100001" ,
        218 => "111100001" ,
        219 => "111100001" ,
        220 => "111100001" ,
        221 => "111100000" ,
        222 => "111100000" ,
        223 => "111100000" ,
        224 => "111100000" ,
        225 => "111100000" ,
        226 => "111100000" ,
        227 => "111100000" ,
        228 => "111011111" ,
        229 => "111011111" ,
        230 => "111011111" ,
        231 => "111011111" ,
        232 => "111011111" ,
        233 => "111011111" ,
        234 => "111011111" ,
        235 => "111011110" ,
        236 => "111011110" ,
        237 => "111011110" ,
        238 => "111011110" ,
        239 => "111011110" ,
        240 => "111011110" ,
        241 => "111011110" ,
        242 => "111011101" ,
        243 => "111011101" ,
        244 => "111011101" ,
        245 => "111011101" ,
        246 => "111011101" ,
        247 => "111011101" ,
        248 => "111011101" ,
        249 => "111011100" ,
        250 => "111011100" ,
        251 => "111011100" ,
        252 => "111011100" ,
        253 => "111011100" ,
        254 => "111011100" ,
        255 => "111011100"
    );

begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <= mem(to_integer(unsigned(address))); 
        end if;
    end process rom;

end architecture synth_c9;

