-------------------------------------------------------------------------------
-- Synthesizable syncronous 8-bit in 8-bit out ROM.
-- Outputs the input multiplied by c2 (as an unsigned integer).
-- 
-- Based on code by M. Treseler available at:
-- http://mysite.ncnetwork.net/reszotzl/sync_rom.vhd
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_rom_c2 is
    generic (data_length : natural := 8;
             add_length  : natural := 8);

    port ( clk          : in  std_logic;
           address      : in  std_logic_vector(add_length-1 downto 0);
           data_out     : out std_logic_vector(data_length-1 downto 0)
       );
end sync_rom_c2;

architecture synth_c2 of sync_rom_c2 is ---------------------------------------------
    constant mem_size : natural := 2**add_length;
    type     mem_type is array (mem_size-1 downto 0) of
    std_logic_vector (data_length-1 downto 0);
    constant mem : mem_type := (
        0 => "00000000" ,
        1 => "00000001" ,
        2 => "00000001" ,
        3 => "00000010" ,
        4 => "00000010" ,
        5 => "00000011" ,
        6 => "00000011" ,
        7 => "00000100" ,
        8 => "00000100" ,
        9 => "00000101" ,
        10 => "00000101" ,
        11 => "00000110" ,
        12 => "00000110" ,
        13 => "00000111" ,
        14 => "00000111" ,
        15 => "00001000" ,
        16 => "00001000" ,
        17 => "00001001" ,
        18 => "00001001" ,
        19 => "00001010" ,
        20 => "00001010" ,
        21 => "00001011" ,
        22 => "00001011" ,
        23 => "00001100" ,
        24 => "00001100" ,
        25 => "00001101" ,
        26 => "00001101" ,
        27 => "00001110" ,
        28 => "00001110" ,
        29 => "00001111" ,
        30 => "00001111" ,
        31 => "00010000" ,
        32 => "00010000" ,
        33 => "00010001" ,
        34 => "00010001" ,
        35 => "00010010" ,
        36 => "00010010" ,
        37 => "00010011" ,
        38 => "00010011" ,
        39 => "00010100" ,
        40 => "00010100" ,
        41 => "00010101" ,
        42 => "00010101" ,
        43 => "00010110" ,
        44 => "00010110" ,
        45 => "00010111" ,
        46 => "00010111" ,
        47 => "00011000" ,
        48 => "00011000" ,
        49 => "00011001" ,
        50 => "00011001" ,
        51 => "00011010" ,
        52 => "00011010" ,
        53 => "00011011" ,
        54 => "00011011" ,
        55 => "00011100" ,
        56 => "00011100" ,
        57 => "00011101" ,
        58 => "00011101" ,
        59 => "00011110" ,
        60 => "00011110" ,
        61 => "00011111" ,
        62 => "00011111" ,
        63 => "00100000" ,
        64 => "00100000" ,
        65 => "00100001" ,
        66 => "00100001" ,
        67 => "00100010" ,
        68 => "00100010" ,
        69 => "00100011" ,
        70 => "00100011" ,
        71 => "00100100" ,
        72 => "00100100" ,
        73 => "00100101" ,
        74 => "00100101" ,
        75 => "00100110" ,
        76 => "00100110" ,
        77 => "00100111" ,
        78 => "00100111" ,
        79 => "00101000" ,
        80 => "00101000" ,
        81 => "00101001" ,
        82 => "00101001" ,
        83 => "00101010" ,
        84 => "00101010" ,
        85 => "00101011" ,
        86 => "00101011" ,
        87 => "00101100" ,
        88 => "00101100" ,
        89 => "00101101" ,
        90 => "00101101" ,
        91 => "00101110" ,
        92 => "00101110" ,
        93 => "00101111" ,
        94 => "00101111" ,
        95 => "00110000" ,
        96 => "00110000" ,
        97 => "00110001" ,
        98 => "00110001" ,
        99 => "00110010" ,
        100 => "00110010" ,
        101 => "00110011" ,
        102 => "00110011" ,
        103 => "00110100" ,
        104 => "00110100" ,
        105 => "00110101" ,
        106 => "00110101" ,
        107 => "00110110" ,
        108 => "00110110" ,
        109 => "00110111" ,
        110 => "00110111" ,
        111 => "00111000" ,
        112 => "00111000" ,
        113 => "00111001" ,
        114 => "00111001" ,
        115 => "00111010" ,
        116 => "00111010" ,
        117 => "00111011" ,
        118 => "00111011" ,
        119 => "00111100" ,
        120 => "00111100" ,
        121 => "00111101" ,
        122 => "00111110" ,
        123 => "00111110" ,
        124 => "00111111" ,
        125 => "00111111" ,
        126 => "01000000" ,
        127 => "01000000" ,
        128 => "01000001" ,
        129 => "01000001" ,
        130 => "01000010" ,
        131 => "01000010" ,
        132 => "01000011" ,
        133 => "01000011" ,
        134 => "01000100" ,
        135 => "01000100" ,
        136 => "01000101" ,
        137 => "01000101" ,
        138 => "01000110" ,
        139 => "01000110" ,
        140 => "01000111" ,
        141 => "01000111" ,
        142 => "01001000" ,
        143 => "01001000" ,
        144 => "01001001" ,
        145 => "01001001" ,
        146 => "01001010" ,
        147 => "01001010" ,
        148 => "01001011" ,
        149 => "01001011" ,
        150 => "01001100" ,
        151 => "01001100" ,
        152 => "01001101" ,
        153 => "01001101" ,
        154 => "01001110" ,
        155 => "01001110" ,
        156 => "01001111" ,
        157 => "01001111" ,
        158 => "01010000" ,
        159 => "01010000" ,
        160 => "01010001" ,
        161 => "01010001" ,
        162 => "01010010" ,
        163 => "01010010" ,
        164 => "01010011" ,
        165 => "01010011" ,
        166 => "01010100" ,
        167 => "01010100" ,
        168 => "01010101" ,
        169 => "01010101" ,
        170 => "01010110" ,
        171 => "01010110" ,
        172 => "01010111" ,
        173 => "01010111" ,
        174 => "01011000" ,
        175 => "01011000" ,
        176 => "01011001" ,
        177 => "01011001" ,
        178 => "01011010" ,
        179 => "01011010" ,
        180 => "01011011" ,
        181 => "01011011" ,
        182 => "01011100" ,
        183 => "01011100" ,
        184 => "01011101" ,
        185 => "01011101" ,
        186 => "01011110" ,
        187 => "01011110" ,
        188 => "01011111" ,
        189 => "01011111" ,
        190 => "01100000" ,
        191 => "01100000" ,
        192 => "01100001" ,
        193 => "01100001" ,
        194 => "01100010" ,
        195 => "01100010" ,
        196 => "01100011" ,
        197 => "01100011" ,
        198 => "01100100" ,
        199 => "01100100" ,
        200 => "01100101" ,
        201 => "01100101" ,
        202 => "01100110" ,
        203 => "01100110" ,
        204 => "01100111" ,
        205 => "01100111" ,
        206 => "01101000" ,
        207 => "01101000" ,
        208 => "01101001" ,
        209 => "01101001" ,
        210 => "01101010" ,
        211 => "01101010" ,
        212 => "01101011" ,
        213 => "01101011" ,
        214 => "01101100" ,
        215 => "01101100" ,
        216 => "01101101" ,
        217 => "01101101" ,
        218 => "01101110" ,
        219 => "01101110" ,
        220 => "01101111" ,
        221 => "01101111" ,
        222 => "01110000" ,
        223 => "01110000" ,
        224 => "01110001" ,
        225 => "01110001" ,
        226 => "01110010" ,
        227 => "01110010" ,
        228 => "01110011" ,
        229 => "01110011" ,
        230 => "01110100" ,
        231 => "01110100" ,
        232 => "01110101" ,
        233 => "01110101" ,
        234 => "01110110" ,
        235 => "01110110" ,
        236 => "01110111" ,
        237 => "01110111" ,
        238 => "01111000" ,
        239 => "01111000" ,
        240 => "01111001" ,
        241 => "01111001" ,
        242 => "01111010" ,
        243 => "01111011" ,
        244 => "01111011" ,
        245 => "01111100" ,
        246 => "01111100" ,
        247 => "01111101" ,
        248 => "01111101" ,
        249 => "01111110" ,
        250 => "01111110" ,
        251 => "01111111" ,
        252 => "01111111" ,
        253 => "10000000" ,
        254 => "10000000" ,
        255 => "10000001"
    );

begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <= mem(to_integer(unsigned(address))); 
        end if;
    end process rom;

end architecture synth_c2;

